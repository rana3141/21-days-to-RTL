// Design and verify mux